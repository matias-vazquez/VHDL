library ieee;
use ieee.std_logic_1164.all;

entity gumnut_system is
  port ( clk_i : in std_logic;
         rst_i : in std_logic );  -- add ports for I/O
end entity gumnut_system;
